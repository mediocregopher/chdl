ENTITY CHIP9684 IS
    PORT(SIGNAL_IN9685 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9686 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9687 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9688 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9689 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9690 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9691 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9692 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9693 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9684;

ARCHITECTURE ARCH OF CHIP9684 IS
    SIGNAL SIGNAL9694 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9694 <= SIGNAL_IN9688;
    SIGNAL_OUT9693 <= SIGNAL_IN9687;
    SIGNAL_OUT9692 <= SIGNAL_IN9686;
    SIGNAL_OUT9691 <= (SIGNAL_IN9686 + ((((SIGNAL_IN9685 + ((SIGNAL_IN9686 and SIGNAL_IN9687) or ((not SIGNAL_IN9686) and SIGNAL_IN9688))) + TO_UNSIGNED(3614090360, 32)) + SIGNAL_IN9689) rol 7));
    SIGNAL9694 <= SIGNAL_IN9688;
END ARCHITECTURE ARCH;


ENTITY CHIP9695 IS
    PORT(SIGNAL_IN9696 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9697 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9698 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9699 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9700 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9701 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9702 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9703 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9704 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9695;

ARCHITECTURE ARCH OF CHIP9695 IS
    SIGNAL SIGNAL9705 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9705 <= SIGNAL_IN9699;
    SIGNAL_OUT9704 <= SIGNAL_IN9698;
    SIGNAL_OUT9703 <= SIGNAL_IN9697;
    SIGNAL_OUT9702 <= (SIGNAL_IN9697 + ((((SIGNAL_IN9696 + ((SIGNAL_IN9697 and SIGNAL_IN9698) or ((not SIGNAL_IN9697) and SIGNAL_IN9699))) + TO_UNSIGNED(3905402710, 32)) + SIGNAL_IN9700) rol 12));
    SIGNAL9705 <= SIGNAL_IN9699;
END ARCHITECTURE ARCH;


ENTITY CHIP9706 IS
    PORT(SIGNAL_IN9707 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9708 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9709 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9710 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9711 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9712 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9713 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9714 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9715 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9706;

ARCHITECTURE ARCH OF CHIP9706 IS
    SIGNAL SIGNAL9716 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9716 <= SIGNAL_IN9710;
    SIGNAL_OUT9715 <= SIGNAL_IN9709;
    SIGNAL_OUT9714 <= SIGNAL_IN9708;
    SIGNAL_OUT9713 <= (SIGNAL_IN9708 + ((((SIGNAL_IN9707 + ((SIGNAL_IN9708 and SIGNAL_IN9709) or ((not SIGNAL_IN9708) and SIGNAL_IN9710))) + TO_UNSIGNED(606105819, 32)) + SIGNAL_IN9711) rol 17));
    SIGNAL9716 <= SIGNAL_IN9710;
END ARCHITECTURE ARCH;


ENTITY CHIP9717 IS
    PORT(SIGNAL_IN9718 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9719 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9720 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9721 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9722 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9723 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9724 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9725 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9726 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9717;

ARCHITECTURE ARCH OF CHIP9717 IS
    SIGNAL SIGNAL9727 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9727 <= SIGNAL_IN9721;
    SIGNAL_OUT9726 <= SIGNAL_IN9720;
    SIGNAL_OUT9725 <= SIGNAL_IN9719;
    SIGNAL_OUT9724 <= (SIGNAL_IN9719 + ((((SIGNAL_IN9718 + ((SIGNAL_IN9719 and SIGNAL_IN9720) or ((not SIGNAL_IN9719) and SIGNAL_IN9721))) + TO_UNSIGNED(3250441966, 32)) + SIGNAL_IN9722) rol 22));
    SIGNAL9727 <= SIGNAL_IN9721;
END ARCHITECTURE ARCH;


ENTITY CHIP9728 IS
    PORT(SIGNAL_IN9729 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9730 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9731 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9732 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9733 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9734 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9735 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9736 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9737 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9728;

ARCHITECTURE ARCH OF CHIP9728 IS
    SIGNAL SIGNAL9738 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9738 <= SIGNAL_IN9732;
    SIGNAL_OUT9737 <= SIGNAL_IN9731;
    SIGNAL_OUT9736 <= SIGNAL_IN9730;
    SIGNAL_OUT9735 <= (SIGNAL_IN9730 + ((((SIGNAL_IN9729 + ((SIGNAL_IN9730 and SIGNAL_IN9731) or ((not SIGNAL_IN9730) and SIGNAL_IN9732))) + TO_UNSIGNED(4118548399, 32)) + SIGNAL_IN9733) rol 7));
    SIGNAL9738 <= SIGNAL_IN9732;
END ARCHITECTURE ARCH;


ENTITY CHIP9739 IS
    PORT(SIGNAL_IN9740 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9741 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9742 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9743 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9744 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9745 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9746 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9747 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9748 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9739;

ARCHITECTURE ARCH OF CHIP9739 IS
    SIGNAL SIGNAL9749 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9749 <= SIGNAL_IN9743;
    SIGNAL_OUT9748 <= SIGNAL_IN9742;
    SIGNAL_OUT9747 <= SIGNAL_IN9741;
    SIGNAL_OUT9746 <= (SIGNAL_IN9741 + ((((SIGNAL_IN9740 + ((SIGNAL_IN9741 and SIGNAL_IN9742) or ((not SIGNAL_IN9741) and SIGNAL_IN9743))) + TO_UNSIGNED(1200080426, 32)) + SIGNAL_IN9744) rol 12));
    SIGNAL9749 <= SIGNAL_IN9743;
END ARCHITECTURE ARCH;


ENTITY CHIP9750 IS
    PORT(SIGNAL_IN9751 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9752 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9753 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9754 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9755 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9756 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9757 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9758 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9759 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9750;

ARCHITECTURE ARCH OF CHIP9750 IS
    SIGNAL SIGNAL9760 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9760 <= SIGNAL_IN9754;
    SIGNAL_OUT9759 <= SIGNAL_IN9753;
    SIGNAL_OUT9758 <= SIGNAL_IN9752;
    SIGNAL_OUT9757 <= (SIGNAL_IN9752 + ((((SIGNAL_IN9751 + ((SIGNAL_IN9752 and SIGNAL_IN9753) or ((not SIGNAL_IN9752) and SIGNAL_IN9754))) + TO_UNSIGNED(2821735955, 32)) + SIGNAL_IN9755) rol 17));
    SIGNAL9760 <= SIGNAL_IN9754;
END ARCHITECTURE ARCH;


ENTITY CHIP9761 IS
    PORT(SIGNAL_IN9762 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9763 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9764 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9765 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9766 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9767 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9768 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9769 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9770 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9761;

ARCHITECTURE ARCH OF CHIP9761 IS
    SIGNAL SIGNAL9771 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9771 <= SIGNAL_IN9765;
    SIGNAL_OUT9770 <= SIGNAL_IN9764;
    SIGNAL_OUT9769 <= SIGNAL_IN9763;
    SIGNAL_OUT9768 <= (SIGNAL_IN9763 + ((((SIGNAL_IN9762 + ((SIGNAL_IN9763 and SIGNAL_IN9764) or ((not SIGNAL_IN9763) and SIGNAL_IN9765))) + TO_UNSIGNED(4249261313, 32)) + SIGNAL_IN9766) rol 22));
    SIGNAL9771 <= SIGNAL_IN9765;
END ARCHITECTURE ARCH;


ENTITY CHIP9772 IS
    PORT(SIGNAL_IN9773 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9774 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9775 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9776 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9777 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9778 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9779 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9780 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9781 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9772;

ARCHITECTURE ARCH OF CHIP9772 IS
    SIGNAL SIGNAL9782 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9782 <= SIGNAL_IN9776;
    SIGNAL_OUT9781 <= SIGNAL_IN9775;
    SIGNAL_OUT9780 <= SIGNAL_IN9774;
    SIGNAL_OUT9779 <= (SIGNAL_IN9774 + ((((SIGNAL_IN9773 + ((SIGNAL_IN9774 and SIGNAL_IN9775) or ((not SIGNAL_IN9774) and SIGNAL_IN9776))) + TO_UNSIGNED(1770035416, 32)) + SIGNAL_IN9777) rol 7));
    SIGNAL9782 <= SIGNAL_IN9776;
END ARCHITECTURE ARCH;


ENTITY CHIP9783 IS
    PORT(SIGNAL_IN9784 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9785 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9786 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9787 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9788 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9789 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9790 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9791 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9792 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9783;

ARCHITECTURE ARCH OF CHIP9783 IS
    SIGNAL SIGNAL9793 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9793 <= SIGNAL_IN9787;
    SIGNAL_OUT9792 <= SIGNAL_IN9786;
    SIGNAL_OUT9791 <= SIGNAL_IN9785;
    SIGNAL_OUT9790 <= (SIGNAL_IN9785 + ((((SIGNAL_IN9784 + ((SIGNAL_IN9785 and SIGNAL_IN9786) or ((not SIGNAL_IN9785) and SIGNAL_IN9787))) + TO_UNSIGNED(2336552879, 32)) + SIGNAL_IN9788) rol 12));
    SIGNAL9793 <= SIGNAL_IN9787;
END ARCHITECTURE ARCH;


ENTITY CHIP9794 IS
    PORT(SIGNAL_IN9795 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9796 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9797 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9798 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9799 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9800 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9801 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9802 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9803 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9794;

ARCHITECTURE ARCH OF CHIP9794 IS
    SIGNAL SIGNAL9804 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9804 <= SIGNAL_IN9798;
    SIGNAL_OUT9803 <= SIGNAL_IN9797;
    SIGNAL_OUT9802 <= SIGNAL_IN9796;
    SIGNAL_OUT9801 <= (SIGNAL_IN9796 + ((((SIGNAL_IN9795 + ((SIGNAL_IN9796 and SIGNAL_IN9797) or ((not SIGNAL_IN9796) and SIGNAL_IN9798))) + TO_UNSIGNED(4294925233, 32)) + SIGNAL_IN9799) rol 17));
    SIGNAL9804 <= SIGNAL_IN9798;
END ARCHITECTURE ARCH;


ENTITY CHIP9805 IS
    PORT(SIGNAL_IN9806 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9807 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9808 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9809 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9810 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9811 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9812 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9813 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9814 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9805;

ARCHITECTURE ARCH OF CHIP9805 IS
    SIGNAL SIGNAL9815 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9815 <= SIGNAL_IN9809;
    SIGNAL_OUT9814 <= SIGNAL_IN9808;
    SIGNAL_OUT9813 <= SIGNAL_IN9807;
    SIGNAL_OUT9812 <= (SIGNAL_IN9807 + ((((SIGNAL_IN9806 + ((SIGNAL_IN9807 and SIGNAL_IN9808) or ((not SIGNAL_IN9807) and SIGNAL_IN9809))) + TO_UNSIGNED(2304563134, 32)) + SIGNAL_IN9810) rol 22));
    SIGNAL9815 <= SIGNAL_IN9809;
END ARCHITECTURE ARCH;


ENTITY CHIP9816 IS
    PORT(SIGNAL_IN9817 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9818 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9819 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9820 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9821 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9822 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9823 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9824 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9825 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9816;

ARCHITECTURE ARCH OF CHIP9816 IS
    SIGNAL SIGNAL9826 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9826 <= SIGNAL_IN9820;
    SIGNAL_OUT9825 <= SIGNAL_IN9819;
    SIGNAL_OUT9824 <= SIGNAL_IN9818;
    SIGNAL_OUT9823 <= (SIGNAL_IN9818 + ((((SIGNAL_IN9817 + ((SIGNAL_IN9818 and SIGNAL_IN9819) or ((not SIGNAL_IN9818) and SIGNAL_IN9820))) + TO_UNSIGNED(1804603682, 32)) + SIGNAL_IN9821) rol 7));
    SIGNAL9826 <= SIGNAL_IN9820;
END ARCHITECTURE ARCH;


ENTITY CHIP9827 IS
    PORT(SIGNAL_IN9828 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9829 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9830 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9831 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9832 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9833 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9834 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9835 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9836 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9827;

ARCHITECTURE ARCH OF CHIP9827 IS
    SIGNAL SIGNAL9837 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9837 <= SIGNAL_IN9831;
    SIGNAL_OUT9836 <= SIGNAL_IN9830;
    SIGNAL_OUT9835 <= SIGNAL_IN9829;
    SIGNAL_OUT9834 <= (SIGNAL_IN9829 + ((((SIGNAL_IN9828 + ((SIGNAL_IN9829 and SIGNAL_IN9830) or ((not SIGNAL_IN9829) and SIGNAL_IN9831))) + TO_UNSIGNED(4254626195, 32)) + SIGNAL_IN9832) rol 12));
    SIGNAL9837 <= SIGNAL_IN9831;
END ARCHITECTURE ARCH;


ENTITY CHIP9838 IS
    PORT(SIGNAL_IN9839 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9840 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9841 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9842 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9843 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9844 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9845 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9846 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9847 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9838;

ARCHITECTURE ARCH OF CHIP9838 IS
    SIGNAL SIGNAL9848 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9848 <= SIGNAL_IN9842;
    SIGNAL_OUT9847 <= SIGNAL_IN9841;
    SIGNAL_OUT9846 <= SIGNAL_IN9840;
    SIGNAL_OUT9845 <= (SIGNAL_IN9840 + ((((SIGNAL_IN9839 + ((SIGNAL_IN9840 and SIGNAL_IN9841) or ((not SIGNAL_IN9840) and SIGNAL_IN9842))) + TO_UNSIGNED(2792965006, 32)) + SIGNAL_IN9843) rol 17));
    SIGNAL9848 <= SIGNAL_IN9842;
END ARCHITECTURE ARCH;


ENTITY CHIP9849 IS
    PORT(SIGNAL_IN9850 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9851 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9852 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9853 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9854 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9855 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9856 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9857 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9858 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9849;

ARCHITECTURE ARCH OF CHIP9849 IS
    SIGNAL SIGNAL9859 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9859 <= SIGNAL_IN9853;
    SIGNAL_OUT9858 <= SIGNAL_IN9852;
    SIGNAL_OUT9857 <= SIGNAL_IN9851;
    SIGNAL_OUT9856 <= (SIGNAL_IN9851 + ((((SIGNAL_IN9850 + ((SIGNAL_IN9851 and SIGNAL_IN9852) or ((not SIGNAL_IN9851) and SIGNAL_IN9853))) + TO_UNSIGNED(1236535329, 32)) + SIGNAL_IN9854) rol 22));
    SIGNAL9859 <= SIGNAL_IN9853;
END ARCHITECTURE ARCH;


ENTITY CHIP9860 IS
    PORT(SIGNAL_IN9861 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9862 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9863 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9864 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9865 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9866 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9867 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9868 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9869 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9860;

ARCHITECTURE ARCH OF CHIP9860 IS
    SIGNAL SIGNAL9870 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9870 <= SIGNAL_IN9864;
    SIGNAL_OUT9869 <= SIGNAL_IN9863;
    SIGNAL_OUT9868 <= SIGNAL_IN9862;
    SIGNAL_OUT9867 <= (SIGNAL_IN9862 + ((((SIGNAL_IN9861 + ((SIGNAL_IN9864 and SIGNAL_IN9862) or ((not SIGNAL_IN9864) and SIGNAL_IN9863))) + TO_UNSIGNED(4129170786, 32)) + SIGNAL_IN9865) rol 5));
    SIGNAL9870 <= SIGNAL_IN9864;
END ARCHITECTURE ARCH;


ENTITY CHIP9871 IS
    PORT(SIGNAL_IN9872 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9873 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9874 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9875 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9876 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9877 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9878 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9879 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9880 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9871;

ARCHITECTURE ARCH OF CHIP9871 IS
    SIGNAL SIGNAL9881 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9881 <= SIGNAL_IN9875;
    SIGNAL_OUT9880 <= SIGNAL_IN9874;
    SIGNAL_OUT9879 <= SIGNAL_IN9873;
    SIGNAL_OUT9878 <= (SIGNAL_IN9873 + ((((SIGNAL_IN9872 + ((SIGNAL_IN9875 and SIGNAL_IN9873) or ((not SIGNAL_IN9875) and SIGNAL_IN9874))) + TO_UNSIGNED(3225465664, 32)) + SIGNAL_IN9876) rol 9));
    SIGNAL9881 <= SIGNAL_IN9875;
END ARCHITECTURE ARCH;


ENTITY CHIP9882 IS
    PORT(SIGNAL_IN9883 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9884 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9885 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9886 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9887 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9888 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9889 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9890 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9891 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9882;

ARCHITECTURE ARCH OF CHIP9882 IS
    SIGNAL SIGNAL9892 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9892 <= SIGNAL_IN9886;
    SIGNAL_OUT9891 <= SIGNAL_IN9885;
    SIGNAL_OUT9890 <= SIGNAL_IN9884;
    SIGNAL_OUT9889 <= (SIGNAL_IN9884 + ((((SIGNAL_IN9883 + ((SIGNAL_IN9886 and SIGNAL_IN9884) or ((not SIGNAL_IN9886) and SIGNAL_IN9885))) + TO_UNSIGNED(643717713, 32)) + SIGNAL_IN9887) rol 14));
    SIGNAL9892 <= SIGNAL_IN9886;
END ARCHITECTURE ARCH;


ENTITY CHIP9893 IS
    PORT(SIGNAL_IN9894 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9895 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9896 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9897 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9898 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9899 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9900 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9901 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9902 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9893;

ARCHITECTURE ARCH OF CHIP9893 IS
    SIGNAL SIGNAL9903 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9903 <= SIGNAL_IN9897;
    SIGNAL_OUT9902 <= SIGNAL_IN9896;
    SIGNAL_OUT9901 <= SIGNAL_IN9895;
    SIGNAL_OUT9900 <= (SIGNAL_IN9895 + ((((SIGNAL_IN9894 + ((SIGNAL_IN9897 and SIGNAL_IN9895) or ((not SIGNAL_IN9897) and SIGNAL_IN9896))) + TO_UNSIGNED(3921069994, 32)) + SIGNAL_IN9898) rol 20));
    SIGNAL9903 <= SIGNAL_IN9897;
END ARCHITECTURE ARCH;


ENTITY CHIP9904 IS
    PORT(SIGNAL_IN9905 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9906 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9907 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9908 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9909 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9910 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9911 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9912 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9913 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9904;

ARCHITECTURE ARCH OF CHIP9904 IS
    SIGNAL SIGNAL9914 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9914 <= SIGNAL_IN9908;
    SIGNAL_OUT9913 <= SIGNAL_IN9907;
    SIGNAL_OUT9912 <= SIGNAL_IN9906;
    SIGNAL_OUT9911 <= (SIGNAL_IN9906 + ((((SIGNAL_IN9905 + ((SIGNAL_IN9908 and SIGNAL_IN9906) or ((not SIGNAL_IN9908) and SIGNAL_IN9907))) + TO_UNSIGNED(3593408605, 32)) + SIGNAL_IN9909) rol 5));
    SIGNAL9914 <= SIGNAL_IN9908;
END ARCHITECTURE ARCH;


ENTITY CHIP9915 IS
    PORT(SIGNAL_IN9916 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9917 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9918 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9919 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9920 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9921 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9922 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9923 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9924 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9915;

ARCHITECTURE ARCH OF CHIP9915 IS
    SIGNAL SIGNAL9925 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9925 <= SIGNAL_IN9919;
    SIGNAL_OUT9924 <= SIGNAL_IN9918;
    SIGNAL_OUT9923 <= SIGNAL_IN9917;
    SIGNAL_OUT9922 <= (SIGNAL_IN9917 + ((((SIGNAL_IN9916 + ((SIGNAL_IN9919 and SIGNAL_IN9917) or ((not SIGNAL_IN9919) and SIGNAL_IN9918))) + TO_UNSIGNED(38016083, 32)) + SIGNAL_IN9920) rol 9));
    SIGNAL9925 <= SIGNAL_IN9919;
END ARCHITECTURE ARCH;


ENTITY CHIP9926 IS
    PORT(SIGNAL_IN9927 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9928 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9929 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9930 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9931 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9932 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9933 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9934 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9935 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9926;

ARCHITECTURE ARCH OF CHIP9926 IS
    SIGNAL SIGNAL9936 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9936 <= SIGNAL_IN9930;
    SIGNAL_OUT9935 <= SIGNAL_IN9929;
    SIGNAL_OUT9934 <= SIGNAL_IN9928;
    SIGNAL_OUT9933 <= (SIGNAL_IN9928 + ((((SIGNAL_IN9927 + ((SIGNAL_IN9930 and SIGNAL_IN9928) or ((not SIGNAL_IN9930) and SIGNAL_IN9929))) + TO_UNSIGNED(3634488961, 32)) + SIGNAL_IN9931) rol 14));
    SIGNAL9936 <= SIGNAL_IN9930;
END ARCHITECTURE ARCH;


ENTITY CHIP9937 IS
    PORT(SIGNAL_IN9938 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9939 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9940 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9941 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9942 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9943 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9944 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9945 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9946 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9937;

ARCHITECTURE ARCH OF CHIP9937 IS
    SIGNAL SIGNAL9947 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9947 <= SIGNAL_IN9941;
    SIGNAL_OUT9946 <= SIGNAL_IN9940;
    SIGNAL_OUT9945 <= SIGNAL_IN9939;
    SIGNAL_OUT9944 <= (SIGNAL_IN9939 + ((((SIGNAL_IN9938 + ((SIGNAL_IN9941 and SIGNAL_IN9939) or ((not SIGNAL_IN9941) and SIGNAL_IN9940))) + TO_UNSIGNED(3889429448, 32)) + SIGNAL_IN9942) rol 20));
    SIGNAL9947 <= SIGNAL_IN9941;
END ARCHITECTURE ARCH;


ENTITY CHIP9948 IS
    PORT(SIGNAL_IN9949 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9950 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9951 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9952 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9953 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9954 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9955 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9956 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9957 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9948;

ARCHITECTURE ARCH OF CHIP9948 IS
    SIGNAL SIGNAL9958 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9958 <= SIGNAL_IN9952;
    SIGNAL_OUT9957 <= SIGNAL_IN9951;
    SIGNAL_OUT9956 <= SIGNAL_IN9950;
    SIGNAL_OUT9955 <= (SIGNAL_IN9950 + ((((SIGNAL_IN9949 + ((SIGNAL_IN9952 and SIGNAL_IN9950) or ((not SIGNAL_IN9952) and SIGNAL_IN9951))) + TO_UNSIGNED(568446438, 32)) + SIGNAL_IN9953) rol 5));
    SIGNAL9958 <= SIGNAL_IN9952;
END ARCHITECTURE ARCH;


ENTITY CHIP9959 IS
    PORT(SIGNAL_IN9960 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9961 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9962 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9963 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9964 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9965 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9966 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9967 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9968 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9959;

ARCHITECTURE ARCH OF CHIP9959 IS
    SIGNAL SIGNAL9969 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9969 <= SIGNAL_IN9963;
    SIGNAL_OUT9968 <= SIGNAL_IN9962;
    SIGNAL_OUT9967 <= SIGNAL_IN9961;
    SIGNAL_OUT9966 <= (SIGNAL_IN9961 + ((((SIGNAL_IN9960 + ((SIGNAL_IN9963 and SIGNAL_IN9961) or ((not SIGNAL_IN9963) and SIGNAL_IN9962))) + TO_UNSIGNED(3275163606, 32)) + SIGNAL_IN9964) rol 9));
    SIGNAL9969 <= SIGNAL_IN9963;
END ARCHITECTURE ARCH;


ENTITY CHIP9970 IS
    PORT(SIGNAL_IN9971 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9972 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9973 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9974 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9975 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9976 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9977 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9978 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9979 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9970;

ARCHITECTURE ARCH OF CHIP9970 IS
    SIGNAL SIGNAL9980 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9980 <= SIGNAL_IN9974;
    SIGNAL_OUT9979 <= SIGNAL_IN9973;
    SIGNAL_OUT9978 <= SIGNAL_IN9972;
    SIGNAL_OUT9977 <= (SIGNAL_IN9972 + ((((SIGNAL_IN9971 + ((SIGNAL_IN9974 and SIGNAL_IN9972) or ((not SIGNAL_IN9974) and SIGNAL_IN9973))) + TO_UNSIGNED(4107603335, 32)) + SIGNAL_IN9975) rol 14));
    SIGNAL9980 <= SIGNAL_IN9974;
END ARCHITECTURE ARCH;


ENTITY CHIP9981 IS
    PORT(SIGNAL_IN9982 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9983 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9984 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9985 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9986 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9987 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9988 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9989 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9990 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9981;

ARCHITECTURE ARCH OF CHIP9981 IS
    SIGNAL SIGNAL9991 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9991 <= SIGNAL_IN9985;
    SIGNAL_OUT9990 <= SIGNAL_IN9984;
    SIGNAL_OUT9989 <= SIGNAL_IN9983;
    SIGNAL_OUT9988 <= (SIGNAL_IN9983 + ((((SIGNAL_IN9982 + ((SIGNAL_IN9985 and SIGNAL_IN9983) or ((not SIGNAL_IN9985) and SIGNAL_IN9984))) + TO_UNSIGNED(1163531501, 32)) + SIGNAL_IN9986) rol 20));
    SIGNAL9991 <= SIGNAL_IN9985;
END ARCHITECTURE ARCH;


ENTITY CHIP9992 IS
    PORT(SIGNAL_IN9993 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9994 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9995 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9996 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9997 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT9998 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9999 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10000 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10001 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9992;

ARCHITECTURE ARCH OF CHIP9992 IS
    SIGNAL SIGNAL10002 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10002 <= SIGNAL_IN9996;
    SIGNAL_OUT10001 <= SIGNAL_IN9995;
    SIGNAL_OUT10000 <= SIGNAL_IN9994;
    SIGNAL_OUT9999 <= (SIGNAL_IN9994 + ((((SIGNAL_IN9993 + ((SIGNAL_IN9996 and SIGNAL_IN9994) or ((not SIGNAL_IN9996) and SIGNAL_IN9995))) + TO_UNSIGNED(2850285829, 32)) + SIGNAL_IN9997) rol 5));
    SIGNAL10002 <= SIGNAL_IN9996;
END ARCHITECTURE ARCH;


ENTITY CHIP10003 IS
    PORT(SIGNAL_IN10004 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10005 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10006 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10007 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10008 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10009 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10010 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10011 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10012 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10003;

ARCHITECTURE ARCH OF CHIP10003 IS
    SIGNAL SIGNAL10013 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10013 <= SIGNAL_IN10007;
    SIGNAL_OUT10012 <= SIGNAL_IN10006;
    SIGNAL_OUT10011 <= SIGNAL_IN10005;
    SIGNAL_OUT10010 <= (SIGNAL_IN10005 + ((((SIGNAL_IN10004 + ((SIGNAL_IN10007 and SIGNAL_IN10005) or ((not SIGNAL_IN10007) and SIGNAL_IN10006))) + TO_UNSIGNED(4243563512, 32)) + SIGNAL_IN10008) rol 9));
    SIGNAL10013 <= SIGNAL_IN10007;
END ARCHITECTURE ARCH;


ENTITY CHIP10014 IS
    PORT(SIGNAL_IN10015 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10016 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10017 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10018 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10019 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10020 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10021 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10022 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10023 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10014;

ARCHITECTURE ARCH OF CHIP10014 IS
    SIGNAL SIGNAL10024 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10024 <= SIGNAL_IN10018;
    SIGNAL_OUT10023 <= SIGNAL_IN10017;
    SIGNAL_OUT10022 <= SIGNAL_IN10016;
    SIGNAL_OUT10021 <= (SIGNAL_IN10016 + ((((SIGNAL_IN10015 + ((SIGNAL_IN10018 and SIGNAL_IN10016) or ((not SIGNAL_IN10018) and SIGNAL_IN10017))) + TO_UNSIGNED(1735328473, 32)) + SIGNAL_IN10019) rol 14));
    SIGNAL10024 <= SIGNAL_IN10018;
END ARCHITECTURE ARCH;


ENTITY CHIP10025 IS
    PORT(SIGNAL_IN10026 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10027 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10028 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10029 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10030 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10031 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10032 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10033 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10034 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10025;

ARCHITECTURE ARCH OF CHIP10025 IS
    SIGNAL SIGNAL10035 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10035 <= SIGNAL_IN10029;
    SIGNAL_OUT10034 <= SIGNAL_IN10028;
    SIGNAL_OUT10033 <= SIGNAL_IN10027;
    SIGNAL_OUT10032 <= (SIGNAL_IN10027 + ((((SIGNAL_IN10026 + ((SIGNAL_IN10029 and SIGNAL_IN10027) or ((not SIGNAL_IN10029) and SIGNAL_IN10028))) + TO_UNSIGNED(2368359562, 32)) + SIGNAL_IN10030) rol 20));
    SIGNAL10035 <= SIGNAL_IN10029;
END ARCHITECTURE ARCH;


ENTITY CHIP10036 IS
    PORT(SIGNAL_IN10037 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10038 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10039 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10040 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10041 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10042 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10043 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10044 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10045 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10036;

ARCHITECTURE ARCH OF CHIP10036 IS
    SIGNAL SIGNAL10046 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10046 <= SIGNAL_IN10040;
    SIGNAL_OUT10045 <= SIGNAL_IN10039;
    SIGNAL_OUT10044 <= SIGNAL_IN10038;
    SIGNAL_OUT10043 <= (SIGNAL_IN10038 + ((((SIGNAL_IN10037 + (SIGNAL_IN10038 xor (SIGNAL_IN10039 xor SIGNAL_IN10040))) + TO_UNSIGNED(4294588738, 32)) + SIGNAL_IN10041) rol 4));
    SIGNAL10046 <= SIGNAL_IN10040;
END ARCHITECTURE ARCH;


ENTITY CHIP10047 IS
    PORT(SIGNAL_IN10048 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10049 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10050 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10051 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10052 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10053 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10054 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10055 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10056 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10047;

ARCHITECTURE ARCH OF CHIP10047 IS
    SIGNAL SIGNAL10057 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10057 <= SIGNAL_IN10051;
    SIGNAL_OUT10056 <= SIGNAL_IN10050;
    SIGNAL_OUT10055 <= SIGNAL_IN10049;
    SIGNAL_OUT10054 <= (SIGNAL_IN10049 + ((((SIGNAL_IN10048 + (SIGNAL_IN10049 xor (SIGNAL_IN10050 xor SIGNAL_IN10051))) + TO_UNSIGNED(2272392833, 32)) + SIGNAL_IN10052) rol 11));
    SIGNAL10057 <= SIGNAL_IN10051;
END ARCHITECTURE ARCH;


ENTITY CHIP10058 IS
    PORT(SIGNAL_IN10059 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10060 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10061 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10062 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10063 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10064 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10065 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10066 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10067 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10058;

ARCHITECTURE ARCH OF CHIP10058 IS
    SIGNAL SIGNAL10068 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10068 <= SIGNAL_IN10062;
    SIGNAL_OUT10067 <= SIGNAL_IN10061;
    SIGNAL_OUT10066 <= SIGNAL_IN10060;
    SIGNAL_OUT10065 <= (SIGNAL_IN10060 + ((((SIGNAL_IN10059 + (SIGNAL_IN10060 xor (SIGNAL_IN10061 xor SIGNAL_IN10062))) + TO_UNSIGNED(1839030562, 32)) + SIGNAL_IN10063) rol 16));
    SIGNAL10068 <= SIGNAL_IN10062;
END ARCHITECTURE ARCH;


ENTITY CHIP10069 IS
    PORT(SIGNAL_IN10070 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10071 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10072 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10073 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10074 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10075 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10076 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10077 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10078 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10069;

ARCHITECTURE ARCH OF CHIP10069 IS
    SIGNAL SIGNAL10079 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10079 <= SIGNAL_IN10073;
    SIGNAL_OUT10078 <= SIGNAL_IN10072;
    SIGNAL_OUT10077 <= SIGNAL_IN10071;
    SIGNAL_OUT10076 <= (SIGNAL_IN10071 + ((((SIGNAL_IN10070 + (SIGNAL_IN10071 xor (SIGNAL_IN10072 xor SIGNAL_IN10073))) + TO_UNSIGNED(4259657740, 32)) + SIGNAL_IN10074) rol 23));
    SIGNAL10079 <= SIGNAL_IN10073;
END ARCHITECTURE ARCH;


ENTITY CHIP10080 IS
    PORT(SIGNAL_IN10081 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10082 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10083 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10084 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10085 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10086 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10087 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10088 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10089 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10080;

ARCHITECTURE ARCH OF CHIP10080 IS
    SIGNAL SIGNAL10090 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10090 <= SIGNAL_IN10084;
    SIGNAL_OUT10089 <= SIGNAL_IN10083;
    SIGNAL_OUT10088 <= SIGNAL_IN10082;
    SIGNAL_OUT10087 <= (SIGNAL_IN10082 + ((((SIGNAL_IN10081 + (SIGNAL_IN10082 xor (SIGNAL_IN10083 xor SIGNAL_IN10084))) + TO_UNSIGNED(2763975236, 32)) + SIGNAL_IN10085) rol 4));
    SIGNAL10090 <= SIGNAL_IN10084;
END ARCHITECTURE ARCH;


ENTITY CHIP10091 IS
    PORT(SIGNAL_IN10092 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10093 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10094 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10095 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10096 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10097 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10098 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10099 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10100 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10091;

ARCHITECTURE ARCH OF CHIP10091 IS
    SIGNAL SIGNAL10101 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10101 <= SIGNAL_IN10095;
    SIGNAL_OUT10100 <= SIGNAL_IN10094;
    SIGNAL_OUT10099 <= SIGNAL_IN10093;
    SIGNAL_OUT10098 <= (SIGNAL_IN10093 + ((((SIGNAL_IN10092 + (SIGNAL_IN10093 xor (SIGNAL_IN10094 xor SIGNAL_IN10095))) + TO_UNSIGNED(1272893353, 32)) + SIGNAL_IN10096) rol 11));
    SIGNAL10101 <= SIGNAL_IN10095;
END ARCHITECTURE ARCH;


ENTITY CHIP10102 IS
    PORT(SIGNAL_IN10103 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10104 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10105 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10106 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10107 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10108 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10109 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10110 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10111 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10102;

ARCHITECTURE ARCH OF CHIP10102 IS
    SIGNAL SIGNAL10112 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10112 <= SIGNAL_IN10106;
    SIGNAL_OUT10111 <= SIGNAL_IN10105;
    SIGNAL_OUT10110 <= SIGNAL_IN10104;
    SIGNAL_OUT10109 <= (SIGNAL_IN10104 + ((((SIGNAL_IN10103 + (SIGNAL_IN10104 xor (SIGNAL_IN10105 xor SIGNAL_IN10106))) + TO_UNSIGNED(4139469664, 32)) + SIGNAL_IN10107) rol 16));
    SIGNAL10112 <= SIGNAL_IN10106;
END ARCHITECTURE ARCH;


ENTITY CHIP10113 IS
    PORT(SIGNAL_IN10114 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10115 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10116 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10117 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10118 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10119 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10120 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10121 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10122 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10113;

ARCHITECTURE ARCH OF CHIP10113 IS
    SIGNAL SIGNAL10123 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10123 <= SIGNAL_IN10117;
    SIGNAL_OUT10122 <= SIGNAL_IN10116;
    SIGNAL_OUT10121 <= SIGNAL_IN10115;
    SIGNAL_OUT10120 <= (SIGNAL_IN10115 + ((((SIGNAL_IN10114 + (SIGNAL_IN10115 xor (SIGNAL_IN10116 xor SIGNAL_IN10117))) + TO_UNSIGNED(3200236656, 32)) + SIGNAL_IN10118) rol 23));
    SIGNAL10123 <= SIGNAL_IN10117;
END ARCHITECTURE ARCH;


ENTITY CHIP10124 IS
    PORT(SIGNAL_IN10125 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10126 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10127 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10128 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10129 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10130 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10131 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10132 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10133 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10124;

ARCHITECTURE ARCH OF CHIP10124 IS
    SIGNAL SIGNAL10134 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10134 <= SIGNAL_IN10128;
    SIGNAL_OUT10133 <= SIGNAL_IN10127;
    SIGNAL_OUT10132 <= SIGNAL_IN10126;
    SIGNAL_OUT10131 <= (SIGNAL_IN10126 + ((((SIGNAL_IN10125 + (SIGNAL_IN10126 xor (SIGNAL_IN10127 xor SIGNAL_IN10128))) + TO_UNSIGNED(681279174, 32)) + SIGNAL_IN10129) rol 4));
    SIGNAL10134 <= SIGNAL_IN10128;
END ARCHITECTURE ARCH;


ENTITY CHIP10135 IS
    PORT(SIGNAL_IN10136 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10137 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10138 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10139 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10140 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10141 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10142 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10143 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10144 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10135;

ARCHITECTURE ARCH OF CHIP10135 IS
    SIGNAL SIGNAL10145 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10145 <= SIGNAL_IN10139;
    SIGNAL_OUT10144 <= SIGNAL_IN10138;
    SIGNAL_OUT10143 <= SIGNAL_IN10137;
    SIGNAL_OUT10142 <= (SIGNAL_IN10137 + ((((SIGNAL_IN10136 + (SIGNAL_IN10137 xor (SIGNAL_IN10138 xor SIGNAL_IN10139))) + TO_UNSIGNED(3936430074, 32)) + SIGNAL_IN10140) rol 11));
    SIGNAL10145 <= SIGNAL_IN10139;
END ARCHITECTURE ARCH;


ENTITY CHIP10146 IS
    PORT(SIGNAL_IN10147 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10148 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10149 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10150 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10151 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10152 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10153 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10154 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10155 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10146;

ARCHITECTURE ARCH OF CHIP10146 IS
    SIGNAL SIGNAL10156 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10156 <= SIGNAL_IN10150;
    SIGNAL_OUT10155 <= SIGNAL_IN10149;
    SIGNAL_OUT10154 <= SIGNAL_IN10148;
    SIGNAL_OUT10153 <= (SIGNAL_IN10148 + ((((SIGNAL_IN10147 + (SIGNAL_IN10148 xor (SIGNAL_IN10149 xor SIGNAL_IN10150))) + TO_UNSIGNED(3572445317, 32)) + SIGNAL_IN10151) rol 16));
    SIGNAL10156 <= SIGNAL_IN10150;
END ARCHITECTURE ARCH;


ENTITY CHIP10157 IS
    PORT(SIGNAL_IN10158 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10159 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10160 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10161 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10162 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10163 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10164 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10165 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10166 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10157;

ARCHITECTURE ARCH OF CHIP10157 IS
    SIGNAL SIGNAL10167 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10167 <= SIGNAL_IN10161;
    SIGNAL_OUT10166 <= SIGNAL_IN10160;
    SIGNAL_OUT10165 <= SIGNAL_IN10159;
    SIGNAL_OUT10164 <= (SIGNAL_IN10159 + ((((SIGNAL_IN10158 + (SIGNAL_IN10159 xor (SIGNAL_IN10160 xor SIGNAL_IN10161))) + TO_UNSIGNED(76029189, 32)) + SIGNAL_IN10162) rol 23));
    SIGNAL10167 <= SIGNAL_IN10161;
END ARCHITECTURE ARCH;


ENTITY CHIP10168 IS
    PORT(SIGNAL_IN10169 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10170 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10171 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10172 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10173 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10174 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10175 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10176 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10177 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10168;

ARCHITECTURE ARCH OF CHIP10168 IS
    SIGNAL SIGNAL10178 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10178 <= SIGNAL_IN10172;
    SIGNAL_OUT10177 <= SIGNAL_IN10171;
    SIGNAL_OUT10176 <= SIGNAL_IN10170;
    SIGNAL_OUT10175 <= (SIGNAL_IN10170 + ((((SIGNAL_IN10169 + (SIGNAL_IN10170 xor (SIGNAL_IN10171 xor SIGNAL_IN10172))) + TO_UNSIGNED(3654602809, 32)) + SIGNAL_IN10173) rol 4));
    SIGNAL10178 <= SIGNAL_IN10172;
END ARCHITECTURE ARCH;


ENTITY CHIP10179 IS
    PORT(SIGNAL_IN10180 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10181 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10182 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10183 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10184 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10185 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10186 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10187 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10188 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10179;

ARCHITECTURE ARCH OF CHIP10179 IS
    SIGNAL SIGNAL10189 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10189 <= SIGNAL_IN10183;
    SIGNAL_OUT10188 <= SIGNAL_IN10182;
    SIGNAL_OUT10187 <= SIGNAL_IN10181;
    SIGNAL_OUT10186 <= (SIGNAL_IN10181 + ((((SIGNAL_IN10180 + (SIGNAL_IN10181 xor (SIGNAL_IN10182 xor SIGNAL_IN10183))) + TO_UNSIGNED(3873151461, 32)) + SIGNAL_IN10184) rol 11));
    SIGNAL10189 <= SIGNAL_IN10183;
END ARCHITECTURE ARCH;


ENTITY CHIP10190 IS
    PORT(SIGNAL_IN10191 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10192 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10193 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10194 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10195 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10196 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10197 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10198 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10199 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10190;

ARCHITECTURE ARCH OF CHIP10190 IS
    SIGNAL SIGNAL10200 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10200 <= SIGNAL_IN10194;
    SIGNAL_OUT10199 <= SIGNAL_IN10193;
    SIGNAL_OUT10198 <= SIGNAL_IN10192;
    SIGNAL_OUT10197 <= (SIGNAL_IN10192 + ((((SIGNAL_IN10191 + (SIGNAL_IN10192 xor (SIGNAL_IN10193 xor SIGNAL_IN10194))) + TO_UNSIGNED(530742520, 32)) + SIGNAL_IN10195) rol 16));
    SIGNAL10200 <= SIGNAL_IN10194;
END ARCHITECTURE ARCH;


ENTITY CHIP10201 IS
    PORT(SIGNAL_IN10202 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10203 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10204 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10205 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10206 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10207 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10208 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10209 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10210 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10201;

ARCHITECTURE ARCH OF CHIP10201 IS
    SIGNAL SIGNAL10211 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10211 <= SIGNAL_IN10205;
    SIGNAL_OUT10210 <= SIGNAL_IN10204;
    SIGNAL_OUT10209 <= SIGNAL_IN10203;
    SIGNAL_OUT10208 <= (SIGNAL_IN10203 + ((((SIGNAL_IN10202 + (SIGNAL_IN10203 xor (SIGNAL_IN10204 xor SIGNAL_IN10205))) + TO_UNSIGNED(3299628645, 32)) + SIGNAL_IN10206) rol 23));
    SIGNAL10211 <= SIGNAL_IN10205;
END ARCHITECTURE ARCH;


ENTITY CHIP10212 IS
    PORT(SIGNAL_IN10213 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10214 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10215 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10216 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10217 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10218 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10219 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10220 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10221 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10212;

ARCHITECTURE ARCH OF CHIP10212 IS
    SIGNAL SIGNAL10222 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10222 <= SIGNAL_IN10216;
    SIGNAL_OUT10221 <= SIGNAL_IN10215;
    SIGNAL_OUT10220 <= SIGNAL_IN10214;
    SIGNAL_OUT10219 <= (SIGNAL_IN10214 + ((((SIGNAL_IN10213 + (SIGNAL_IN10215 xor (SIGNAL_IN10214 or (not SIGNAL_IN10216)))) + TO_UNSIGNED(4096336452, 32)) + SIGNAL_IN10217) rol 6));
    SIGNAL10222 <= SIGNAL_IN10216;
END ARCHITECTURE ARCH;


ENTITY CHIP10223 IS
    PORT(SIGNAL_IN10224 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10225 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10226 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10227 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10228 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10229 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10230 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10231 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10232 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10223;

ARCHITECTURE ARCH OF CHIP10223 IS
    SIGNAL SIGNAL10233 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10233 <= SIGNAL_IN10227;
    SIGNAL_OUT10232 <= SIGNAL_IN10226;
    SIGNAL_OUT10231 <= SIGNAL_IN10225;
    SIGNAL_OUT10230 <= (SIGNAL_IN10225 + ((((SIGNAL_IN10224 + (SIGNAL_IN10226 xor (SIGNAL_IN10225 or (not SIGNAL_IN10227)))) + TO_UNSIGNED(1126891415, 32)) + SIGNAL_IN10228) rol 10));
    SIGNAL10233 <= SIGNAL_IN10227;
END ARCHITECTURE ARCH;


ENTITY CHIP10234 IS
    PORT(SIGNAL_IN10235 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10236 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10237 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10238 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10239 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10240 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10241 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10242 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10243 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10234;

ARCHITECTURE ARCH OF CHIP10234 IS
    SIGNAL SIGNAL10244 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10244 <= SIGNAL_IN10238;
    SIGNAL_OUT10243 <= SIGNAL_IN10237;
    SIGNAL_OUT10242 <= SIGNAL_IN10236;
    SIGNAL_OUT10241 <= (SIGNAL_IN10236 + ((((SIGNAL_IN10235 + (SIGNAL_IN10237 xor (SIGNAL_IN10236 or (not SIGNAL_IN10238)))) + TO_UNSIGNED(2878612391, 32)) + SIGNAL_IN10239) rol 15));
    SIGNAL10244 <= SIGNAL_IN10238;
END ARCHITECTURE ARCH;


ENTITY CHIP10245 IS
    PORT(SIGNAL_IN10246 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10247 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10248 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10249 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10250 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10251 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10252 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10253 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10254 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10245;

ARCHITECTURE ARCH OF CHIP10245 IS
    SIGNAL SIGNAL10255 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10255 <= SIGNAL_IN10249;
    SIGNAL_OUT10254 <= SIGNAL_IN10248;
    SIGNAL_OUT10253 <= SIGNAL_IN10247;
    SIGNAL_OUT10252 <= (SIGNAL_IN10247 + ((((SIGNAL_IN10246 + (SIGNAL_IN10248 xor (SIGNAL_IN10247 or (not SIGNAL_IN10249)))) + TO_UNSIGNED(4237533241, 32)) + SIGNAL_IN10250) rol 21));
    SIGNAL10255 <= SIGNAL_IN10249;
END ARCHITECTURE ARCH;


ENTITY CHIP10256 IS
    PORT(SIGNAL_IN10257 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10258 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10259 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10260 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10261 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10262 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10263 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10264 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10265 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10256;

ARCHITECTURE ARCH OF CHIP10256 IS
    SIGNAL SIGNAL10266 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10266 <= SIGNAL_IN10260;
    SIGNAL_OUT10265 <= SIGNAL_IN10259;
    SIGNAL_OUT10264 <= SIGNAL_IN10258;
    SIGNAL_OUT10263 <= (SIGNAL_IN10258 + ((((SIGNAL_IN10257 + (SIGNAL_IN10259 xor (SIGNAL_IN10258 or (not SIGNAL_IN10260)))) + TO_UNSIGNED(1700485571, 32)) + SIGNAL_IN10261) rol 6));
    SIGNAL10266 <= SIGNAL_IN10260;
END ARCHITECTURE ARCH;


ENTITY CHIP10267 IS
    PORT(SIGNAL_IN10268 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10269 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10270 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10271 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10272 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10273 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10274 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10275 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10276 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10267;

ARCHITECTURE ARCH OF CHIP10267 IS
    SIGNAL SIGNAL10277 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10277 <= SIGNAL_IN10271;
    SIGNAL_OUT10276 <= SIGNAL_IN10270;
    SIGNAL_OUT10275 <= SIGNAL_IN10269;
    SIGNAL_OUT10274 <= (SIGNAL_IN10269 + ((((SIGNAL_IN10268 + (SIGNAL_IN10270 xor (SIGNAL_IN10269 or (not SIGNAL_IN10271)))) + TO_UNSIGNED(2399980690, 32)) + SIGNAL_IN10272) rol 10));
    SIGNAL10277 <= SIGNAL_IN10271;
END ARCHITECTURE ARCH;


ENTITY CHIP10278 IS
    PORT(SIGNAL_IN10279 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10280 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10281 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10282 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10283 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10284 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10285 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10286 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10287 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10278;

ARCHITECTURE ARCH OF CHIP10278 IS
    SIGNAL SIGNAL10288 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10288 <= SIGNAL_IN10282;
    SIGNAL_OUT10287 <= SIGNAL_IN10281;
    SIGNAL_OUT10286 <= SIGNAL_IN10280;
    SIGNAL_OUT10285 <= (SIGNAL_IN10280 + ((((SIGNAL_IN10279 + (SIGNAL_IN10281 xor (SIGNAL_IN10280 or (not SIGNAL_IN10282)))) + TO_UNSIGNED(4293915773, 32)) + SIGNAL_IN10283) rol 15));
    SIGNAL10288 <= SIGNAL_IN10282;
END ARCHITECTURE ARCH;


ENTITY CHIP10289 IS
    PORT(SIGNAL_IN10290 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10291 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10292 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10293 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10294 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10295 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10296 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10297 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10298 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10289;

ARCHITECTURE ARCH OF CHIP10289 IS
    SIGNAL SIGNAL10299 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10299 <= SIGNAL_IN10293;
    SIGNAL_OUT10298 <= SIGNAL_IN10292;
    SIGNAL_OUT10297 <= SIGNAL_IN10291;
    SIGNAL_OUT10296 <= (SIGNAL_IN10291 + ((((SIGNAL_IN10290 + (SIGNAL_IN10292 xor (SIGNAL_IN10291 or (not SIGNAL_IN10293)))) + TO_UNSIGNED(2240044497, 32)) + SIGNAL_IN10294) rol 21));
    SIGNAL10299 <= SIGNAL_IN10293;
END ARCHITECTURE ARCH;


ENTITY CHIP10300 IS
    PORT(SIGNAL_IN10301 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10302 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10303 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10304 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10305 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10306 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10307 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10308 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10309 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10300;

ARCHITECTURE ARCH OF CHIP10300 IS
    SIGNAL SIGNAL10310 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10310 <= SIGNAL_IN10304;
    SIGNAL_OUT10309 <= SIGNAL_IN10303;
    SIGNAL_OUT10308 <= SIGNAL_IN10302;
    SIGNAL_OUT10307 <= (SIGNAL_IN10302 + ((((SIGNAL_IN10301 + (SIGNAL_IN10303 xor (SIGNAL_IN10302 or (not SIGNAL_IN10304)))) + TO_UNSIGNED(1873313359, 32)) + SIGNAL_IN10305) rol 6));
    SIGNAL10310 <= SIGNAL_IN10304;
END ARCHITECTURE ARCH;


ENTITY CHIP10311 IS
    PORT(SIGNAL_IN10312 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10313 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10314 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10315 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10316 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10317 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10318 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10319 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10320 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10311;

ARCHITECTURE ARCH OF CHIP10311 IS
    SIGNAL SIGNAL10321 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10321 <= SIGNAL_IN10315;
    SIGNAL_OUT10320 <= SIGNAL_IN10314;
    SIGNAL_OUT10319 <= SIGNAL_IN10313;
    SIGNAL_OUT10318 <= (SIGNAL_IN10313 + ((((SIGNAL_IN10312 + (SIGNAL_IN10314 xor (SIGNAL_IN10313 or (not SIGNAL_IN10315)))) + TO_UNSIGNED(4264355552, 32)) + SIGNAL_IN10316) rol 10));
    SIGNAL10321 <= SIGNAL_IN10315;
END ARCHITECTURE ARCH;


ENTITY CHIP10322 IS
    PORT(SIGNAL_IN10323 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10324 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10325 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10326 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10327 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10328 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10329 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10330 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10331 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10322;

ARCHITECTURE ARCH OF CHIP10322 IS
    SIGNAL SIGNAL10332 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10332 <= SIGNAL_IN10326;
    SIGNAL_OUT10331 <= SIGNAL_IN10325;
    SIGNAL_OUT10330 <= SIGNAL_IN10324;
    SIGNAL_OUT10329 <= (SIGNAL_IN10324 + ((((SIGNAL_IN10323 + (SIGNAL_IN10325 xor (SIGNAL_IN10324 or (not SIGNAL_IN10326)))) + TO_UNSIGNED(2734768916, 32)) + SIGNAL_IN10327) rol 15));
    SIGNAL10332 <= SIGNAL_IN10326;
END ARCHITECTURE ARCH;


ENTITY CHIP10333 IS
    PORT(SIGNAL_IN10334 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10335 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10336 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10337 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10338 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10339 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10340 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10341 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10342 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10333;

ARCHITECTURE ARCH OF CHIP10333 IS
    SIGNAL SIGNAL10343 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10343 <= SIGNAL_IN10337;
    SIGNAL_OUT10342 <= SIGNAL_IN10336;
    SIGNAL_OUT10341 <= SIGNAL_IN10335;
    SIGNAL_OUT10340 <= (SIGNAL_IN10335 + ((((SIGNAL_IN10334 + (SIGNAL_IN10336 xor (SIGNAL_IN10335 or (not SIGNAL_IN10337)))) + TO_UNSIGNED(1309151649, 32)) + SIGNAL_IN10338) rol 21));
    SIGNAL10343 <= SIGNAL_IN10337;
END ARCHITECTURE ARCH;


ENTITY CHIP10344 IS
    PORT(SIGNAL_IN10345 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10346 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10347 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10348 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10349 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10350 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10351 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10352 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10353 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10344;

ARCHITECTURE ARCH OF CHIP10344 IS
    SIGNAL SIGNAL10354 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10354 <= SIGNAL_IN10348;
    SIGNAL_OUT10353 <= SIGNAL_IN10347;
    SIGNAL_OUT10352 <= SIGNAL_IN10346;
    SIGNAL_OUT10351 <= (SIGNAL_IN10346 + ((((SIGNAL_IN10345 + (SIGNAL_IN10347 xor (SIGNAL_IN10346 or (not SIGNAL_IN10348)))) + TO_UNSIGNED(4149444226, 32)) + SIGNAL_IN10349) rol 6));
    SIGNAL10354 <= SIGNAL_IN10348;
END ARCHITECTURE ARCH;


ENTITY CHIP10355 IS
    PORT(SIGNAL_IN10356 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10357 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10358 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10359 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10360 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10361 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10362 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10363 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10364 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10355;

ARCHITECTURE ARCH OF CHIP10355 IS
    SIGNAL SIGNAL10365 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10365 <= SIGNAL_IN10359;
    SIGNAL_OUT10364 <= SIGNAL_IN10358;
    SIGNAL_OUT10363 <= SIGNAL_IN10357;
    SIGNAL_OUT10362 <= (SIGNAL_IN10357 + ((((SIGNAL_IN10356 + (SIGNAL_IN10358 xor (SIGNAL_IN10357 or (not SIGNAL_IN10359)))) + TO_UNSIGNED(3174756917, 32)) + SIGNAL_IN10360) rol 10));
    SIGNAL10365 <= SIGNAL_IN10359;
END ARCHITECTURE ARCH;


ENTITY CHIP10366 IS
    PORT(SIGNAL_IN10367 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10368 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10369 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10370 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10371 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10372 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10373 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10374 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10375 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10366;

ARCHITECTURE ARCH OF CHIP10366 IS
    SIGNAL SIGNAL10376 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10376 <= SIGNAL_IN10370;
    SIGNAL_OUT10375 <= SIGNAL_IN10369;
    SIGNAL_OUT10374 <= SIGNAL_IN10368;
    SIGNAL_OUT10373 <= (SIGNAL_IN10368 + ((((SIGNAL_IN10367 + (SIGNAL_IN10369 xor (SIGNAL_IN10368 or (not SIGNAL_IN10370)))) + TO_UNSIGNED(718787259, 32)) + SIGNAL_IN10371) rol 15));
    SIGNAL10376 <= SIGNAL_IN10370;
END ARCHITECTURE ARCH;


ENTITY CHIP10377 IS
    PORT(SIGNAL_IN10378 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10379 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10380 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10381 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN10382 : IN UNSIGNED(31 downto 0);
    SIGNAL_OUT10383 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10384 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10385 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT10386 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP10377;

ARCHITECTURE ARCH OF CHIP10377 IS
    SIGNAL SIGNAL10387 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL10387 <= SIGNAL_IN10381;
    SIGNAL_OUT10386 <= SIGNAL_IN10380;
    SIGNAL_OUT10385 <= SIGNAL_IN10379;
    SIGNAL_OUT10384 <= (SIGNAL_IN10379 + ((((SIGNAL_IN10378 + (SIGNAL_IN10380 xor (SIGNAL_IN10379 or (not SIGNAL_IN10381)))) + TO_UNSIGNED(3951481745, 32)) + SIGNAL_IN10382) rol 21));
    SIGNAL10387 <= SIGNAL_IN10381;
END ARCHITECTURE ARCH;


ENTITY CHIP9398 IS
    PORT(SIGNAL_IN9399 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9400 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9401 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9402 : IN UNSIGNED(31 downto 0);
    SIGNAL_IN9403 : IN STD_LOGIC_VECTOR(511 DOWNTO 0);
    SIGNAL_OUT9404 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9405 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9406 : OUT UNSIGNED(31 downto 0);
    SIGNAL_OUT9407 : OUT UNSIGNED(31 downto 0));
BEGIN
END ENTITY CHIP9398;

ARCHITECTURE ARCH OF CHIP9398 IS
    SIGNAL SIGNAL9408 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9409 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9410 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9411 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9412 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9413 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9414 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9415 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9416 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9417 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9418 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9419 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9420 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9421 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9422 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9423 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9424 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9425 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9426 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9427 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9428 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9429 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9430 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9431 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9432 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9433 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9434 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9435 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9436 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9437 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9438 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9439 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9440 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9441 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9442 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9443 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9444 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9445 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9446 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9447 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9448 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9449 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9450 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9451 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9452 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9453 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9454 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9455 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9456 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9457 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9458 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9459 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9460 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9461 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9462 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9463 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9464 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9465 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9466 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9467 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9468 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9469 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9470 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9471 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9472 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9473 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9474 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9475 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9476 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9477 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9478 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9479 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9480 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9481 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9482 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9483 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9484 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9485 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9486 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9487 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9488 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9489 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9490 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9491 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9492 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9493 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9494 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9495 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9496 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9497 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9498 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9499 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9500 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9501 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9502 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9503 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9504 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9505 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9506 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9507 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9508 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9509 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9510 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9511 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9512 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9513 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9514 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9515 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9516 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9517 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9518 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9519 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9520 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9521 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9522 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9523 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9524 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9525 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9526 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9527 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9528 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9529 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9530 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9531 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9532 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9533 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9534 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9535 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9536 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9537 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9538 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9539 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9540 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9541 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9542 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9543 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9544 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9545 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9546 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9547 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9548 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9549 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9550 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9551 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9552 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9553 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9554 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9555 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9556 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9557 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9558 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9559 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9560 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9561 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9562 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9563 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9564 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9565 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9566 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9567 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9568 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9569 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9570 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9571 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9572 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9573 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9574 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9575 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9576 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9577 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9578 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9579 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9580 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9581 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9582 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9583 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9584 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9585 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9586 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9587 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9588 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9589 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9590 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9591 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9592 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9593 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9594 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9595 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9596 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9597 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9598 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9599 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9600 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9601 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9602 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9603 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9604 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9605 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9606 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9607 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9608 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9609 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9610 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9611 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9612 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9613 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9614 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9615 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9616 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9617 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9618 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9619 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9620 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9621 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9622 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9623 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9624 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9625 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9626 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9627 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9628 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9629 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9630 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9631 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9632 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9633 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9634 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9635 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9636 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9637 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9638 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9639 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9640 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9641 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9642 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9643 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9644 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9645 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9646 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9647 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9648 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9649 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9650 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9651 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9652 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9653 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9654 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9655 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9656 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9657 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9658 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9659 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9660 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9661 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9662 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9663 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9664 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9665 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9666 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9667 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9668 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9669 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9670 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9671 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9672 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9673 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9674 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9675 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9676 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9677 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9678 : UNSIGNED(31 downto 0);
    SIGNAL SIGNAL9679 : UNSIGNED(31 downto 0);
BEGIN
    SIGNAL9408 <= UNSIGNED(SIGNAL_IN9403(31 DOWNTO 0));
    SIGNAL9409 <= UNSIGNED(SIGNAL_IN9403(63 DOWNTO 32));
    SIGNAL9410 <= UNSIGNED(SIGNAL_IN9403(95 DOWNTO 64));
    SIGNAL9411 <= UNSIGNED(SIGNAL_IN9403(127 DOWNTO 96));
    SIGNAL9412 <= UNSIGNED(SIGNAL_IN9403(159 DOWNTO 128));
    SIGNAL9413 <= UNSIGNED(SIGNAL_IN9403(191 DOWNTO 160));
    SIGNAL9414 <= UNSIGNED(SIGNAL_IN9403(223 DOWNTO 192));
    SIGNAL9415 <= UNSIGNED(SIGNAL_IN9403(255 DOWNTO 224));
    SIGNAL9416 <= UNSIGNED(SIGNAL_IN9403(287 DOWNTO 256));
    SIGNAL9417 <= UNSIGNED(SIGNAL_IN9403(319 DOWNTO 288));
    SIGNAL9418 <= UNSIGNED(SIGNAL_IN9403(351 DOWNTO 320));
    SIGNAL9419 <= UNSIGNED(SIGNAL_IN9403(383 DOWNTO 352));
    SIGNAL9420 <= UNSIGNED(SIGNAL_IN9403(415 DOWNTO 384));
    SIGNAL9421 <= UNSIGNED(SIGNAL_IN9403(447 DOWNTO 416));
    SIGNAL9422 <= UNSIGNED(SIGNAL_IN9403(479 DOWNTO 448));
    SIGNAL9423 <= UNSIGNED(SIGNAL_IN9403(511 DOWNTO 480));
    CHIP_INST10388 : ENTITY CHIP9684(ARCH) PORT MAP(SIGNAL_IN9685 => SIGNAL_IN9399
    , SIGNAL_IN9686 => SIGNAL_IN9400
    , SIGNAL_IN9687 => SIGNAL_IN9401
    , SIGNAL_IN9688 => SIGNAL_IN9402
    , SIGNAL_IN9689 => SIGNAL9408
    , SIGNAL_OUT9690 => SIGNAL9425
    , SIGNAL_OUT9691 => SIGNAL9489
    , SIGNAL_OUT9692 => SIGNAL9553
    , SIGNAL_OUT9693 => SIGNAL9617
    );
    CHIP_INST10389 : ENTITY CHIP9695(ARCH) PORT MAP(SIGNAL_IN9696 => SIGNAL9425
    , SIGNAL_IN9697 => SIGNAL9489
    , SIGNAL_IN9698 => SIGNAL9553
    , SIGNAL_IN9699 => SIGNAL9617
    , SIGNAL_IN9700 => SIGNAL9409
    , SIGNAL_OUT9701 => SIGNAL9426
    , SIGNAL_OUT9702 => SIGNAL9490
    , SIGNAL_OUT9703 => SIGNAL9554
    , SIGNAL_OUT9704 => SIGNAL9618
    );
    CHIP_INST10390 : ENTITY CHIP9706(ARCH) PORT MAP(SIGNAL_IN9707 => SIGNAL9426
    , SIGNAL_IN9708 => SIGNAL9490
    , SIGNAL_IN9709 => SIGNAL9554
    , SIGNAL_IN9710 => SIGNAL9618
    , SIGNAL_IN9711 => SIGNAL9410
    , SIGNAL_OUT9712 => SIGNAL9427
    , SIGNAL_OUT9713 => SIGNAL9491
    , SIGNAL_OUT9714 => SIGNAL9555
    , SIGNAL_OUT9715 => SIGNAL9619
    );
    CHIP_INST10391 : ENTITY CHIP9717(ARCH) PORT MAP(SIGNAL_IN9718 => SIGNAL9427
    , SIGNAL_IN9719 => SIGNAL9491
    , SIGNAL_IN9720 => SIGNAL9555
    , SIGNAL_IN9721 => SIGNAL9619
    , SIGNAL_IN9722 => SIGNAL9411
    , SIGNAL_OUT9723 => SIGNAL9428
    , SIGNAL_OUT9724 => SIGNAL9492
    , SIGNAL_OUT9725 => SIGNAL9556
    , SIGNAL_OUT9726 => SIGNAL9620
    );
    CHIP_INST10392 : ENTITY CHIP9728(ARCH) PORT MAP(SIGNAL_IN9729 => SIGNAL9428
    , SIGNAL_IN9730 => SIGNAL9492
    , SIGNAL_IN9731 => SIGNAL9556
    , SIGNAL_IN9732 => SIGNAL9620
    , SIGNAL_IN9733 => SIGNAL9412
    , SIGNAL_OUT9734 => SIGNAL9429
    , SIGNAL_OUT9735 => SIGNAL9493
    , SIGNAL_OUT9736 => SIGNAL9557
    , SIGNAL_OUT9737 => SIGNAL9621
    );
    CHIP_INST10393 : ENTITY CHIP9739(ARCH) PORT MAP(SIGNAL_IN9740 => SIGNAL9429
    , SIGNAL_IN9741 => SIGNAL9493
    , SIGNAL_IN9742 => SIGNAL9557
    , SIGNAL_IN9743 => SIGNAL9621
    , SIGNAL_IN9744 => SIGNAL9413
    , SIGNAL_OUT9745 => SIGNAL9430
    , SIGNAL_OUT9746 => SIGNAL9494
    , SIGNAL_OUT9747 => SIGNAL9558
    , SIGNAL_OUT9748 => SIGNAL9622
    );
    CHIP_INST10394 : ENTITY CHIP9750(ARCH) PORT MAP(SIGNAL_IN9751 => SIGNAL9430
    , SIGNAL_IN9752 => SIGNAL9494
    , SIGNAL_IN9753 => SIGNAL9558
    , SIGNAL_IN9754 => SIGNAL9622
    , SIGNAL_IN9755 => SIGNAL9414
    , SIGNAL_OUT9756 => SIGNAL9431
    , SIGNAL_OUT9757 => SIGNAL9495
    , SIGNAL_OUT9758 => SIGNAL9559
    , SIGNAL_OUT9759 => SIGNAL9623
    );
    CHIP_INST10395 : ENTITY CHIP9761(ARCH) PORT MAP(SIGNAL_IN9762 => SIGNAL9431
    , SIGNAL_IN9763 => SIGNAL9495
    , SIGNAL_IN9764 => SIGNAL9559
    , SIGNAL_IN9765 => SIGNAL9623
    , SIGNAL_IN9766 => SIGNAL9415
    , SIGNAL_OUT9767 => SIGNAL9432
    , SIGNAL_OUT9768 => SIGNAL9496
    , SIGNAL_OUT9769 => SIGNAL9560
    , SIGNAL_OUT9770 => SIGNAL9624
    );
    CHIP_INST10396 : ENTITY CHIP9772(ARCH) PORT MAP(SIGNAL_IN9773 => SIGNAL9432
    , SIGNAL_IN9774 => SIGNAL9496
    , SIGNAL_IN9775 => SIGNAL9560
    , SIGNAL_IN9776 => SIGNAL9624
    , SIGNAL_IN9777 => SIGNAL9416
    , SIGNAL_OUT9778 => SIGNAL9433
    , SIGNAL_OUT9779 => SIGNAL9497
    , SIGNAL_OUT9780 => SIGNAL9561
    , SIGNAL_OUT9781 => SIGNAL9625
    );
    CHIP_INST10397 : ENTITY CHIP9783(ARCH) PORT MAP(SIGNAL_IN9784 => SIGNAL9433
    , SIGNAL_IN9785 => SIGNAL9497
    , SIGNAL_IN9786 => SIGNAL9561
    , SIGNAL_IN9787 => SIGNAL9625
    , SIGNAL_IN9788 => SIGNAL9417
    , SIGNAL_OUT9789 => SIGNAL9434
    , SIGNAL_OUT9790 => SIGNAL9498
    , SIGNAL_OUT9791 => SIGNAL9562
    , SIGNAL_OUT9792 => SIGNAL9626
    );
    CHIP_INST10398 : ENTITY CHIP9794(ARCH) PORT MAP(SIGNAL_IN9795 => SIGNAL9434
    , SIGNAL_IN9796 => SIGNAL9498
    , SIGNAL_IN9797 => SIGNAL9562
    , SIGNAL_IN9798 => SIGNAL9626
    , SIGNAL_IN9799 => SIGNAL9418
    , SIGNAL_OUT9800 => SIGNAL9435
    , SIGNAL_OUT9801 => SIGNAL9499
    , SIGNAL_OUT9802 => SIGNAL9563
    , SIGNAL_OUT9803 => SIGNAL9627
    );
    CHIP_INST10399 : ENTITY CHIP9805(ARCH) PORT MAP(SIGNAL_IN9806 => SIGNAL9435
    , SIGNAL_IN9807 => SIGNAL9499
    , SIGNAL_IN9808 => SIGNAL9563
    , SIGNAL_IN9809 => SIGNAL9627
    , SIGNAL_IN9810 => SIGNAL9419
    , SIGNAL_OUT9811 => SIGNAL9436
    , SIGNAL_OUT9812 => SIGNAL9500
    , SIGNAL_OUT9813 => SIGNAL9564
    , SIGNAL_OUT9814 => SIGNAL9628
    );
    CHIP_INST10400 : ENTITY CHIP9816(ARCH) PORT MAP(SIGNAL_IN9817 => SIGNAL9436
    , SIGNAL_IN9818 => SIGNAL9500
    , SIGNAL_IN9819 => SIGNAL9564
    , SIGNAL_IN9820 => SIGNAL9628
    , SIGNAL_IN9821 => SIGNAL9420
    , SIGNAL_OUT9822 => SIGNAL9437
    , SIGNAL_OUT9823 => SIGNAL9501
    , SIGNAL_OUT9824 => SIGNAL9565
    , SIGNAL_OUT9825 => SIGNAL9629
    );
    CHIP_INST10401 : ENTITY CHIP9827(ARCH) PORT MAP(SIGNAL_IN9828 => SIGNAL9437
    , SIGNAL_IN9829 => SIGNAL9501
    , SIGNAL_IN9830 => SIGNAL9565
    , SIGNAL_IN9831 => SIGNAL9629
    , SIGNAL_IN9832 => SIGNAL9421
    , SIGNAL_OUT9833 => SIGNAL9438
    , SIGNAL_OUT9834 => SIGNAL9502
    , SIGNAL_OUT9835 => SIGNAL9566
    , SIGNAL_OUT9836 => SIGNAL9630
    );
    CHIP_INST10402 : ENTITY CHIP9838(ARCH) PORT MAP(SIGNAL_IN9839 => SIGNAL9438
    , SIGNAL_IN9840 => SIGNAL9502
    , SIGNAL_IN9841 => SIGNAL9566
    , SIGNAL_IN9842 => SIGNAL9630
    , SIGNAL_IN9843 => SIGNAL9422
    , SIGNAL_OUT9844 => SIGNAL9439
    , SIGNAL_OUT9845 => SIGNAL9503
    , SIGNAL_OUT9846 => SIGNAL9567
    , SIGNAL_OUT9847 => SIGNAL9631
    );
    CHIP_INST10403 : ENTITY CHIP9849(ARCH) PORT MAP(SIGNAL_IN9850 => SIGNAL9439
    , SIGNAL_IN9851 => SIGNAL9503
    , SIGNAL_IN9852 => SIGNAL9567
    , SIGNAL_IN9853 => SIGNAL9631
    , SIGNAL_IN9854 => SIGNAL9423
    , SIGNAL_OUT9855 => SIGNAL9440
    , SIGNAL_OUT9856 => SIGNAL9504
    , SIGNAL_OUT9857 => SIGNAL9568
    , SIGNAL_OUT9858 => SIGNAL9632
    );
    CHIP_INST10404 : ENTITY CHIP9860(ARCH) PORT MAP(SIGNAL_IN9861 => SIGNAL9440
    , SIGNAL_IN9862 => SIGNAL9504
    , SIGNAL_IN9863 => SIGNAL9568
    , SIGNAL_IN9864 => SIGNAL9632
    , SIGNAL_IN9865 => SIGNAL9409
    , SIGNAL_OUT9866 => SIGNAL9441
    , SIGNAL_OUT9867 => SIGNAL9505
    , SIGNAL_OUT9868 => SIGNAL9569
    , SIGNAL_OUT9869 => SIGNAL9633
    );
    CHIP_INST10405 : ENTITY CHIP9871(ARCH) PORT MAP(SIGNAL_IN9872 => SIGNAL9441
    , SIGNAL_IN9873 => SIGNAL9505
    , SIGNAL_IN9874 => SIGNAL9569
    , SIGNAL_IN9875 => SIGNAL9633
    , SIGNAL_IN9876 => SIGNAL9414
    , SIGNAL_OUT9877 => SIGNAL9442
    , SIGNAL_OUT9878 => SIGNAL9506
    , SIGNAL_OUT9879 => SIGNAL9570
    , SIGNAL_OUT9880 => SIGNAL9634
    );
    CHIP_INST10406 : ENTITY CHIP9882(ARCH) PORT MAP(SIGNAL_IN9883 => SIGNAL9442
    , SIGNAL_IN9884 => SIGNAL9506
    , SIGNAL_IN9885 => SIGNAL9570
    , SIGNAL_IN9886 => SIGNAL9634
    , SIGNAL_IN9887 => SIGNAL9419
    , SIGNAL_OUT9888 => SIGNAL9443
    , SIGNAL_OUT9889 => SIGNAL9507
    , SIGNAL_OUT9890 => SIGNAL9571
    , SIGNAL_OUT9891 => SIGNAL9635
    );
    CHIP_INST10407 : ENTITY CHIP9893(ARCH) PORT MAP(SIGNAL_IN9894 => SIGNAL9443
    , SIGNAL_IN9895 => SIGNAL9507
    , SIGNAL_IN9896 => SIGNAL9571
    , SIGNAL_IN9897 => SIGNAL9635
    , SIGNAL_IN9898 => SIGNAL9408
    , SIGNAL_OUT9899 => SIGNAL9444
    , SIGNAL_OUT9900 => SIGNAL9508
    , SIGNAL_OUT9901 => SIGNAL9572
    , SIGNAL_OUT9902 => SIGNAL9636
    );
    CHIP_INST10408 : ENTITY CHIP9904(ARCH) PORT MAP(SIGNAL_IN9905 => SIGNAL9444
    , SIGNAL_IN9906 => SIGNAL9508
    , SIGNAL_IN9907 => SIGNAL9572
    , SIGNAL_IN9908 => SIGNAL9636
    , SIGNAL_IN9909 => SIGNAL9413
    , SIGNAL_OUT9910 => SIGNAL9445
    , SIGNAL_OUT9911 => SIGNAL9509
    , SIGNAL_OUT9912 => SIGNAL9573
    , SIGNAL_OUT9913 => SIGNAL9637
    );
    CHIP_INST10409 : ENTITY CHIP9915(ARCH) PORT MAP(SIGNAL_IN9916 => SIGNAL9445
    , SIGNAL_IN9917 => SIGNAL9509
    , SIGNAL_IN9918 => SIGNAL9573
    , SIGNAL_IN9919 => SIGNAL9637
    , SIGNAL_IN9920 => SIGNAL9418
    , SIGNAL_OUT9921 => SIGNAL9446
    , SIGNAL_OUT9922 => SIGNAL9510
    , SIGNAL_OUT9923 => SIGNAL9574
    , SIGNAL_OUT9924 => SIGNAL9638
    );
    CHIP_INST10410 : ENTITY CHIP9926(ARCH) PORT MAP(SIGNAL_IN9927 => SIGNAL9446
    , SIGNAL_IN9928 => SIGNAL9510
    , SIGNAL_IN9929 => SIGNAL9574
    , SIGNAL_IN9930 => SIGNAL9638
    , SIGNAL_IN9931 => SIGNAL9423
    , SIGNAL_OUT9932 => SIGNAL9447
    , SIGNAL_OUT9933 => SIGNAL9511
    , SIGNAL_OUT9934 => SIGNAL9575
    , SIGNAL_OUT9935 => SIGNAL9639
    );
    CHIP_INST10411 : ENTITY CHIP9937(ARCH) PORT MAP(SIGNAL_IN9938 => SIGNAL9447
    , SIGNAL_IN9939 => SIGNAL9511
    , SIGNAL_IN9940 => SIGNAL9575
    , SIGNAL_IN9941 => SIGNAL9639
    , SIGNAL_IN9942 => SIGNAL9412
    , SIGNAL_OUT9943 => SIGNAL9448
    , SIGNAL_OUT9944 => SIGNAL9512
    , SIGNAL_OUT9945 => SIGNAL9576
    , SIGNAL_OUT9946 => SIGNAL9640
    );
    CHIP_INST10412 : ENTITY CHIP9948(ARCH) PORT MAP(SIGNAL_IN9949 => SIGNAL9448
    , SIGNAL_IN9950 => SIGNAL9512
    , SIGNAL_IN9951 => SIGNAL9576
    , SIGNAL_IN9952 => SIGNAL9640
    , SIGNAL_IN9953 => SIGNAL9417
    , SIGNAL_OUT9954 => SIGNAL9449
    , SIGNAL_OUT9955 => SIGNAL9513
    , SIGNAL_OUT9956 => SIGNAL9577
    , SIGNAL_OUT9957 => SIGNAL9641
    );
    CHIP_INST10413 : ENTITY CHIP9959(ARCH) PORT MAP(SIGNAL_IN9960 => SIGNAL9449
    , SIGNAL_IN9961 => SIGNAL9513
    , SIGNAL_IN9962 => SIGNAL9577
    , SIGNAL_IN9963 => SIGNAL9641
    , SIGNAL_IN9964 => SIGNAL9422
    , SIGNAL_OUT9965 => SIGNAL9450
    , SIGNAL_OUT9966 => SIGNAL9514
    , SIGNAL_OUT9967 => SIGNAL9578
    , SIGNAL_OUT9968 => SIGNAL9642
    );
    CHIP_INST10414 : ENTITY CHIP9970(ARCH) PORT MAP(SIGNAL_IN9971 => SIGNAL9450
    , SIGNAL_IN9972 => SIGNAL9514
    , SIGNAL_IN9973 => SIGNAL9578
    , SIGNAL_IN9974 => SIGNAL9642
    , SIGNAL_IN9975 => SIGNAL9411
    , SIGNAL_OUT9976 => SIGNAL9451
    , SIGNAL_OUT9977 => SIGNAL9515
    , SIGNAL_OUT9978 => SIGNAL9579
    , SIGNAL_OUT9979 => SIGNAL9643
    );
    CHIP_INST10415 : ENTITY CHIP9981(ARCH) PORT MAP(SIGNAL_IN9982 => SIGNAL9451
    , SIGNAL_IN9983 => SIGNAL9515
    , SIGNAL_IN9984 => SIGNAL9579
    , SIGNAL_IN9985 => SIGNAL9643
    , SIGNAL_IN9986 => SIGNAL9416
    , SIGNAL_OUT9987 => SIGNAL9452
    , SIGNAL_OUT9988 => SIGNAL9516
    , SIGNAL_OUT9989 => SIGNAL9580
    , SIGNAL_OUT9990 => SIGNAL9644
    );
    CHIP_INST10416 : ENTITY CHIP9992(ARCH) PORT MAP(SIGNAL_IN9993 => SIGNAL9452
    , SIGNAL_IN9994 => SIGNAL9516
    , SIGNAL_IN9995 => SIGNAL9580
    , SIGNAL_IN9996 => SIGNAL9644
    , SIGNAL_IN9997 => SIGNAL9421
    , SIGNAL_OUT9998 => SIGNAL9453
    , SIGNAL_OUT9999 => SIGNAL9517
    , SIGNAL_OUT10000 => SIGNAL9581
    , SIGNAL_OUT10001 => SIGNAL9645
    );
    CHIP_INST10417 : ENTITY CHIP10003(ARCH) PORT MAP(SIGNAL_IN10004 => SIGNAL9453
    , SIGNAL_IN10005 => SIGNAL9517
    , SIGNAL_IN10006 => SIGNAL9581
    , SIGNAL_IN10007 => SIGNAL9645
    , SIGNAL_IN10008 => SIGNAL9410
    , SIGNAL_OUT10009 => SIGNAL9454
    , SIGNAL_OUT10010 => SIGNAL9518
    , SIGNAL_OUT10011 => SIGNAL9582
    , SIGNAL_OUT10012 => SIGNAL9646
    );
    CHIP_INST10418 : ENTITY CHIP10014(ARCH) PORT MAP(SIGNAL_IN10015 => SIGNAL9454
    , SIGNAL_IN10016 => SIGNAL9518
    , SIGNAL_IN10017 => SIGNAL9582
    , SIGNAL_IN10018 => SIGNAL9646
    , SIGNAL_IN10019 => SIGNAL9415
    , SIGNAL_OUT10020 => SIGNAL9455
    , SIGNAL_OUT10021 => SIGNAL9519
    , SIGNAL_OUT10022 => SIGNAL9583
    , SIGNAL_OUT10023 => SIGNAL9647
    );
    CHIP_INST10419 : ENTITY CHIP10025(ARCH) PORT MAP(SIGNAL_IN10026 => SIGNAL9455
    , SIGNAL_IN10027 => SIGNAL9519
    , SIGNAL_IN10028 => SIGNAL9583
    , SIGNAL_IN10029 => SIGNAL9647
    , SIGNAL_IN10030 => SIGNAL9420
    , SIGNAL_OUT10031 => SIGNAL9456
    , SIGNAL_OUT10032 => SIGNAL9520
    , SIGNAL_OUT10033 => SIGNAL9584
    , SIGNAL_OUT10034 => SIGNAL9648
    );
    CHIP_INST10420 : ENTITY CHIP10036(ARCH) PORT MAP(SIGNAL_IN10037 => SIGNAL9456
    , SIGNAL_IN10038 => SIGNAL9520
    , SIGNAL_IN10039 => SIGNAL9584
    , SIGNAL_IN10040 => SIGNAL9648
    , SIGNAL_IN10041 => SIGNAL9413
    , SIGNAL_OUT10042 => SIGNAL9457
    , SIGNAL_OUT10043 => SIGNAL9521
    , SIGNAL_OUT10044 => SIGNAL9585
    , SIGNAL_OUT10045 => SIGNAL9649
    );
    CHIP_INST10421 : ENTITY CHIP10047(ARCH) PORT MAP(SIGNAL_IN10048 => SIGNAL9457
    , SIGNAL_IN10049 => SIGNAL9521
    , SIGNAL_IN10050 => SIGNAL9585
    , SIGNAL_IN10051 => SIGNAL9649
    , SIGNAL_IN10052 => SIGNAL9416
    , SIGNAL_OUT10053 => SIGNAL9458
    , SIGNAL_OUT10054 => SIGNAL9522
    , SIGNAL_OUT10055 => SIGNAL9586
    , SIGNAL_OUT10056 => SIGNAL9650
    );
    CHIP_INST10422 : ENTITY CHIP10058(ARCH) PORT MAP(SIGNAL_IN10059 => SIGNAL9458
    , SIGNAL_IN10060 => SIGNAL9522
    , SIGNAL_IN10061 => SIGNAL9586
    , SIGNAL_IN10062 => SIGNAL9650
    , SIGNAL_IN10063 => SIGNAL9419
    , SIGNAL_OUT10064 => SIGNAL9459
    , SIGNAL_OUT10065 => SIGNAL9523
    , SIGNAL_OUT10066 => SIGNAL9587
    , SIGNAL_OUT10067 => SIGNAL9651
    );
    CHIP_INST10423 : ENTITY CHIP10069(ARCH) PORT MAP(SIGNAL_IN10070 => SIGNAL9459
    , SIGNAL_IN10071 => SIGNAL9523
    , SIGNAL_IN10072 => SIGNAL9587
    , SIGNAL_IN10073 => SIGNAL9651
    , SIGNAL_IN10074 => SIGNAL9422
    , SIGNAL_OUT10075 => SIGNAL9460
    , SIGNAL_OUT10076 => SIGNAL9524
    , SIGNAL_OUT10077 => SIGNAL9588
    , SIGNAL_OUT10078 => SIGNAL9652
    );
    CHIP_INST10424 : ENTITY CHIP10080(ARCH) PORT MAP(SIGNAL_IN10081 => SIGNAL9460
    , SIGNAL_IN10082 => SIGNAL9524
    , SIGNAL_IN10083 => SIGNAL9588
    , SIGNAL_IN10084 => SIGNAL9652
    , SIGNAL_IN10085 => SIGNAL9409
    , SIGNAL_OUT10086 => SIGNAL9461
    , SIGNAL_OUT10087 => SIGNAL9525
    , SIGNAL_OUT10088 => SIGNAL9589
    , SIGNAL_OUT10089 => SIGNAL9653
    );
    CHIP_INST10425 : ENTITY CHIP10091(ARCH) PORT MAP(SIGNAL_IN10092 => SIGNAL9461
    , SIGNAL_IN10093 => SIGNAL9525
    , SIGNAL_IN10094 => SIGNAL9589
    , SIGNAL_IN10095 => SIGNAL9653
    , SIGNAL_IN10096 => SIGNAL9412
    , SIGNAL_OUT10097 => SIGNAL9462
    , SIGNAL_OUT10098 => SIGNAL9526
    , SIGNAL_OUT10099 => SIGNAL9590
    , SIGNAL_OUT10100 => SIGNAL9654
    );
    CHIP_INST10426 : ENTITY CHIP10102(ARCH) PORT MAP(SIGNAL_IN10103 => SIGNAL9462
    , SIGNAL_IN10104 => SIGNAL9526
    , SIGNAL_IN10105 => SIGNAL9590
    , SIGNAL_IN10106 => SIGNAL9654
    , SIGNAL_IN10107 => SIGNAL9415
    , SIGNAL_OUT10108 => SIGNAL9463
    , SIGNAL_OUT10109 => SIGNAL9527
    , SIGNAL_OUT10110 => SIGNAL9591
    , SIGNAL_OUT10111 => SIGNAL9655
    );
    CHIP_INST10427 : ENTITY CHIP10113(ARCH) PORT MAP(SIGNAL_IN10114 => SIGNAL9463
    , SIGNAL_IN10115 => SIGNAL9527
    , SIGNAL_IN10116 => SIGNAL9591
    , SIGNAL_IN10117 => SIGNAL9655
    , SIGNAL_IN10118 => SIGNAL9418
    , SIGNAL_OUT10119 => SIGNAL9464
    , SIGNAL_OUT10120 => SIGNAL9528
    , SIGNAL_OUT10121 => SIGNAL9592
    , SIGNAL_OUT10122 => SIGNAL9656
    );
    CHIP_INST10428 : ENTITY CHIP10124(ARCH) PORT MAP(SIGNAL_IN10125 => SIGNAL9464
    , SIGNAL_IN10126 => SIGNAL9528
    , SIGNAL_IN10127 => SIGNAL9592
    , SIGNAL_IN10128 => SIGNAL9656
    , SIGNAL_IN10129 => SIGNAL9421
    , SIGNAL_OUT10130 => SIGNAL9465
    , SIGNAL_OUT10131 => SIGNAL9529
    , SIGNAL_OUT10132 => SIGNAL9593
    , SIGNAL_OUT10133 => SIGNAL9657
    );
    CHIP_INST10429 : ENTITY CHIP10135(ARCH) PORT MAP(SIGNAL_IN10136 => SIGNAL9465
    , SIGNAL_IN10137 => SIGNAL9529
    , SIGNAL_IN10138 => SIGNAL9593
    , SIGNAL_IN10139 => SIGNAL9657
    , SIGNAL_IN10140 => SIGNAL9408
    , SIGNAL_OUT10141 => SIGNAL9466
    , SIGNAL_OUT10142 => SIGNAL9530
    , SIGNAL_OUT10143 => SIGNAL9594
    , SIGNAL_OUT10144 => SIGNAL9658
    );
    CHIP_INST10430 : ENTITY CHIP10146(ARCH) PORT MAP(SIGNAL_IN10147 => SIGNAL9466
    , SIGNAL_IN10148 => SIGNAL9530
    , SIGNAL_IN10149 => SIGNAL9594
    , SIGNAL_IN10150 => SIGNAL9658
    , SIGNAL_IN10151 => SIGNAL9411
    , SIGNAL_OUT10152 => SIGNAL9467
    , SIGNAL_OUT10153 => SIGNAL9531
    , SIGNAL_OUT10154 => SIGNAL9595
    , SIGNAL_OUT10155 => SIGNAL9659
    );
    CHIP_INST10431 : ENTITY CHIP10157(ARCH) PORT MAP(SIGNAL_IN10158 => SIGNAL9467
    , SIGNAL_IN10159 => SIGNAL9531
    , SIGNAL_IN10160 => SIGNAL9595
    , SIGNAL_IN10161 => SIGNAL9659
    , SIGNAL_IN10162 => SIGNAL9414
    , SIGNAL_OUT10163 => SIGNAL9468
    , SIGNAL_OUT10164 => SIGNAL9532
    , SIGNAL_OUT10165 => SIGNAL9596
    , SIGNAL_OUT10166 => SIGNAL9660
    );
    CHIP_INST10432 : ENTITY CHIP10168(ARCH) PORT MAP(SIGNAL_IN10169 => SIGNAL9468
    , SIGNAL_IN10170 => SIGNAL9532
    , SIGNAL_IN10171 => SIGNAL9596
    , SIGNAL_IN10172 => SIGNAL9660
    , SIGNAL_IN10173 => SIGNAL9417
    , SIGNAL_OUT10174 => SIGNAL9469
    , SIGNAL_OUT10175 => SIGNAL9533
    , SIGNAL_OUT10176 => SIGNAL9597
    , SIGNAL_OUT10177 => SIGNAL9661
    );
    CHIP_INST10433 : ENTITY CHIP10179(ARCH) PORT MAP(SIGNAL_IN10180 => SIGNAL9469
    , SIGNAL_IN10181 => SIGNAL9533
    , SIGNAL_IN10182 => SIGNAL9597
    , SIGNAL_IN10183 => SIGNAL9661
    , SIGNAL_IN10184 => SIGNAL9420
    , SIGNAL_OUT10185 => SIGNAL9470
    , SIGNAL_OUT10186 => SIGNAL9534
    , SIGNAL_OUT10187 => SIGNAL9598
    , SIGNAL_OUT10188 => SIGNAL9662
    );
    CHIP_INST10434 : ENTITY CHIP10190(ARCH) PORT MAP(SIGNAL_IN10191 => SIGNAL9470
    , SIGNAL_IN10192 => SIGNAL9534
    , SIGNAL_IN10193 => SIGNAL9598
    , SIGNAL_IN10194 => SIGNAL9662
    , SIGNAL_IN10195 => SIGNAL9423
    , SIGNAL_OUT10196 => SIGNAL9471
    , SIGNAL_OUT10197 => SIGNAL9535
    , SIGNAL_OUT10198 => SIGNAL9599
    , SIGNAL_OUT10199 => SIGNAL9663
    );
    CHIP_INST10435 : ENTITY CHIP10201(ARCH) PORT MAP(SIGNAL_IN10202 => SIGNAL9471
    , SIGNAL_IN10203 => SIGNAL9535
    , SIGNAL_IN10204 => SIGNAL9599
    , SIGNAL_IN10205 => SIGNAL9663
    , SIGNAL_IN10206 => SIGNAL9410
    , SIGNAL_OUT10207 => SIGNAL9472
    , SIGNAL_OUT10208 => SIGNAL9536
    , SIGNAL_OUT10209 => SIGNAL9600
    , SIGNAL_OUT10210 => SIGNAL9664
    );
    CHIP_INST10436 : ENTITY CHIP10212(ARCH) PORT MAP(SIGNAL_IN10213 => SIGNAL9472
    , SIGNAL_IN10214 => SIGNAL9536
    , SIGNAL_IN10215 => SIGNAL9600
    , SIGNAL_IN10216 => SIGNAL9664
    , SIGNAL_IN10217 => SIGNAL9408
    , SIGNAL_OUT10218 => SIGNAL9473
    , SIGNAL_OUT10219 => SIGNAL9537
    , SIGNAL_OUT10220 => SIGNAL9601
    , SIGNAL_OUT10221 => SIGNAL9665
    );
    CHIP_INST10437 : ENTITY CHIP10223(ARCH) PORT MAP(SIGNAL_IN10224 => SIGNAL9473
    , SIGNAL_IN10225 => SIGNAL9537
    , SIGNAL_IN10226 => SIGNAL9601
    , SIGNAL_IN10227 => SIGNAL9665
    , SIGNAL_IN10228 => SIGNAL9415
    , SIGNAL_OUT10229 => SIGNAL9474
    , SIGNAL_OUT10230 => SIGNAL9538
    , SIGNAL_OUT10231 => SIGNAL9602
    , SIGNAL_OUT10232 => SIGNAL9666
    );
    CHIP_INST10438 : ENTITY CHIP10234(ARCH) PORT MAP(SIGNAL_IN10235 => SIGNAL9474
    , SIGNAL_IN10236 => SIGNAL9538
    , SIGNAL_IN10237 => SIGNAL9602
    , SIGNAL_IN10238 => SIGNAL9666
    , SIGNAL_IN10239 => SIGNAL9422
    , SIGNAL_OUT10240 => SIGNAL9475
    , SIGNAL_OUT10241 => SIGNAL9539
    , SIGNAL_OUT10242 => SIGNAL9603
    , SIGNAL_OUT10243 => SIGNAL9667
    );
    CHIP_INST10439 : ENTITY CHIP10245(ARCH) PORT MAP(SIGNAL_IN10246 => SIGNAL9475
    , SIGNAL_IN10247 => SIGNAL9539
    , SIGNAL_IN10248 => SIGNAL9603
    , SIGNAL_IN10249 => SIGNAL9667
    , SIGNAL_IN10250 => SIGNAL9413
    , SIGNAL_OUT10251 => SIGNAL9476
    , SIGNAL_OUT10252 => SIGNAL9540
    , SIGNAL_OUT10253 => SIGNAL9604
    , SIGNAL_OUT10254 => SIGNAL9668
    );
    CHIP_INST10440 : ENTITY CHIP10256(ARCH) PORT MAP(SIGNAL_IN10257 => SIGNAL9476
    , SIGNAL_IN10258 => SIGNAL9540
    , SIGNAL_IN10259 => SIGNAL9604
    , SIGNAL_IN10260 => SIGNAL9668
    , SIGNAL_IN10261 => SIGNAL9420
    , SIGNAL_OUT10262 => SIGNAL9477
    , SIGNAL_OUT10263 => SIGNAL9541
    , SIGNAL_OUT10264 => SIGNAL9605
    , SIGNAL_OUT10265 => SIGNAL9669
    );
    CHIP_INST10441 : ENTITY CHIP10267(ARCH) PORT MAP(SIGNAL_IN10268 => SIGNAL9477
    , SIGNAL_IN10269 => SIGNAL9541
    , SIGNAL_IN10270 => SIGNAL9605
    , SIGNAL_IN10271 => SIGNAL9669
    , SIGNAL_IN10272 => SIGNAL9411
    , SIGNAL_OUT10273 => SIGNAL9478
    , SIGNAL_OUT10274 => SIGNAL9542
    , SIGNAL_OUT10275 => SIGNAL9606
    , SIGNAL_OUT10276 => SIGNAL9670
    );
    CHIP_INST10442 : ENTITY CHIP10278(ARCH) PORT MAP(SIGNAL_IN10279 => SIGNAL9478
    , SIGNAL_IN10280 => SIGNAL9542
    , SIGNAL_IN10281 => SIGNAL9606
    , SIGNAL_IN10282 => SIGNAL9670
    , SIGNAL_IN10283 => SIGNAL9418
    , SIGNAL_OUT10284 => SIGNAL9479
    , SIGNAL_OUT10285 => SIGNAL9543
    , SIGNAL_OUT10286 => SIGNAL9607
    , SIGNAL_OUT10287 => SIGNAL9671
    );
    CHIP_INST10443 : ENTITY CHIP10289(ARCH) PORT MAP(SIGNAL_IN10290 => SIGNAL9479
    , SIGNAL_IN10291 => SIGNAL9543
    , SIGNAL_IN10292 => SIGNAL9607
    , SIGNAL_IN10293 => SIGNAL9671
    , SIGNAL_IN10294 => SIGNAL9409
    , SIGNAL_OUT10295 => SIGNAL9480
    , SIGNAL_OUT10296 => SIGNAL9544
    , SIGNAL_OUT10297 => SIGNAL9608
    , SIGNAL_OUT10298 => SIGNAL9672
    );
    CHIP_INST10444 : ENTITY CHIP10300(ARCH) PORT MAP(SIGNAL_IN10301 => SIGNAL9480
    , SIGNAL_IN10302 => SIGNAL9544
    , SIGNAL_IN10303 => SIGNAL9608
    , SIGNAL_IN10304 => SIGNAL9672
    , SIGNAL_IN10305 => SIGNAL9416
    , SIGNAL_OUT10306 => SIGNAL9481
    , SIGNAL_OUT10307 => SIGNAL9545
    , SIGNAL_OUT10308 => SIGNAL9609
    , SIGNAL_OUT10309 => SIGNAL9673
    );
    CHIP_INST10445 : ENTITY CHIP10311(ARCH) PORT MAP(SIGNAL_IN10312 => SIGNAL9481
    , SIGNAL_IN10313 => SIGNAL9545
    , SIGNAL_IN10314 => SIGNAL9609
    , SIGNAL_IN10315 => SIGNAL9673
    , SIGNAL_IN10316 => SIGNAL9423
    , SIGNAL_OUT10317 => SIGNAL9482
    , SIGNAL_OUT10318 => SIGNAL9546
    , SIGNAL_OUT10319 => SIGNAL9610
    , SIGNAL_OUT10320 => SIGNAL9674
    );
    CHIP_INST10446 : ENTITY CHIP10322(ARCH) PORT MAP(SIGNAL_IN10323 => SIGNAL9482
    , SIGNAL_IN10324 => SIGNAL9546
    , SIGNAL_IN10325 => SIGNAL9610
    , SIGNAL_IN10326 => SIGNAL9674
    , SIGNAL_IN10327 => SIGNAL9414
    , SIGNAL_OUT10328 => SIGNAL9483
    , SIGNAL_OUT10329 => SIGNAL9547
    , SIGNAL_OUT10330 => SIGNAL9611
    , SIGNAL_OUT10331 => SIGNAL9675
    );
    CHIP_INST10447 : ENTITY CHIP10333(ARCH) PORT MAP(SIGNAL_IN10334 => SIGNAL9483
    , SIGNAL_IN10335 => SIGNAL9547
    , SIGNAL_IN10336 => SIGNAL9611
    , SIGNAL_IN10337 => SIGNAL9675
    , SIGNAL_IN10338 => SIGNAL9421
    , SIGNAL_OUT10339 => SIGNAL9484
    , SIGNAL_OUT10340 => SIGNAL9548
    , SIGNAL_OUT10341 => SIGNAL9612
    , SIGNAL_OUT10342 => SIGNAL9676
    );
    CHIP_INST10448 : ENTITY CHIP10344(ARCH) PORT MAP(SIGNAL_IN10345 => SIGNAL9484
    , SIGNAL_IN10346 => SIGNAL9548
    , SIGNAL_IN10347 => SIGNAL9612
    , SIGNAL_IN10348 => SIGNAL9676
    , SIGNAL_IN10349 => SIGNAL9412
    , SIGNAL_OUT10350 => SIGNAL9485
    , SIGNAL_OUT10351 => SIGNAL9549
    , SIGNAL_OUT10352 => SIGNAL9613
    , SIGNAL_OUT10353 => SIGNAL9677
    );
    CHIP_INST10449 : ENTITY CHIP10355(ARCH) PORT MAP(SIGNAL_IN10356 => SIGNAL9485
    , SIGNAL_IN10357 => SIGNAL9549
    , SIGNAL_IN10358 => SIGNAL9613
    , SIGNAL_IN10359 => SIGNAL9677
    , SIGNAL_IN10360 => SIGNAL9419
    , SIGNAL_OUT10361 => SIGNAL9486
    , SIGNAL_OUT10362 => SIGNAL9550
    , SIGNAL_OUT10363 => SIGNAL9614
    , SIGNAL_OUT10364 => SIGNAL9678
    );
    CHIP_INST10450 : ENTITY CHIP10366(ARCH) PORT MAP(SIGNAL_IN10367 => SIGNAL9486
    , SIGNAL_IN10368 => SIGNAL9550
    , SIGNAL_IN10369 => SIGNAL9614
    , SIGNAL_IN10370 => SIGNAL9678
    , SIGNAL_IN10371 => SIGNAL9410
    , SIGNAL_OUT10372 => SIGNAL9487
    , SIGNAL_OUT10373 => SIGNAL9551
    , SIGNAL_OUT10374 => SIGNAL9615
    , SIGNAL_OUT10375 => SIGNAL9679
    );
    CHIP_INST10451 : ENTITY CHIP10377(ARCH) PORT MAP(SIGNAL_IN10378 => SIGNAL9487
    , SIGNAL_IN10379 => SIGNAL9551
    , SIGNAL_IN10380 => SIGNAL9615
    , SIGNAL_IN10381 => SIGNAL9679
    , SIGNAL_IN10382 => SIGNAL9417
    , SIGNAL_OUT10383 => SIGNAL_OUT9404
    , SIGNAL_OUT10384 => SIGNAL_OUT9405
    , SIGNAL_OUT10385 => SIGNAL_OUT9406
    , SIGNAL_OUT10386 => SIGNAL_OUT9407
    );
END ARCHITECTURE ARCH;

